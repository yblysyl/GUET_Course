LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ADDR IS
PORT(
    I15,I14,I13,I12:IN STD_LOGIC;
    CF,ZF,SF,T4,P1,P2,P3:IN STD_LOGIC;
    SE5,SE4,SE3,SE2,SE1,SE0:OUT STD_LOGIC
);
END ADDR;
ARCHITECTURE A OF ADDR IS 
BEGIN 
    SE5<=NOT((P3 AND ZF AND T4) OR (P3 AND NOT(SF) AND T4));
    SE4<=NOT(P2 AND NOT(ZF) AND T4);
    SE3<=NOT(P1 AND I15 AND T4);
    SE2<=NOT(P1 AND I14 AND T4);
    SE1<=NOT(P1 AND I13 AND T4);
    SE0<=NOT(P1 AND I12 AND T4);
END A;

