LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ROM IS
PORT(
    DOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    ADDR:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    CS_I:IN STD_LOGIC
);
END ROM;
ARCHITECTURE A OF ROM IS
BEGIN
    DOUT<="0010000000000000" WHEN ADDR="00000000" AND CS_I='0' ELSE		--MOV	R0,00H
          "0010000100000101" WHEN ADDR="00000001" AND CS_I='0' ELSE		--MOV	R1,05H
          "0001001000000000" WHEN ADDR="00000010" AND CS_I='0' ELSE		--INPUT:IN1	R2
          "0011100000000000" WHEN ADDR="00000011" AND CS_I='0' ELSE		--STO1	R2,(R0)
          "0100000000000000" WHEN ADDR="00000100" AND CS_I='0' ELSE		--INC		R0
          "0101000100000000" WHEN ADDR="00000101" AND CS_I='0' ELSE		--DEC		R1
          "0110000100000000" WHEN ADDR="00000110" AND CS_I='0' ELSE		--TEST		R1
          "1000000000000010" WHEN ADDR="00000111" AND CS_I='0' ELSE		--JNZ	INPUT
          "0010000000000000" WHEN ADDR="00001000" AND CS_I='0' ELSE		--MOV	R0,00H
          "0010000100000101" WHEN ADDR="00001001" AND CS_I='0' ELSE		--MOV	R1,05H
          "1001001100000000" WHEN ADDR="00001010" AND CS_I='0' ELSE		--LAD (R0),R3
          "1001001000000000" WHEN ADDR="00001011" AND CS_I='0' ELSE		--JUDGE:LAD  (R0),R2
          "0110001000000000" WHEN ADDR="00001100" AND CS_I='0' ELSE		--TEST		R2 
          "1010000000010001" WHEN ADDR="00001101" AND CS_I='0' ELSE		--JNS		YES 
          "0111111000000000" WHEN ADDR="00001110" AND CS_I='0' ELSE		--CMP	R3,R2 
          "1010000000010001" WHEN ADDR="00001111" AND CS_I='0' ELSE		--JNS		YES 
          "1101101100000000" WHEN ADDR="00010000" AND CS_I='0' ELSE		--MOV1  R2,R3 
          "0100000000000000" WHEN ADDR="00010001" AND CS_I='0' ELSE		--YES:INC	R0
          "0101000100000000" WHEN ADDR="00010010" AND CS_I='0' ELSE		--DEC		R1
          "0110000100000000" WHEN ADDR="00010011" AND CS_I='0' ELSE		--TEST		R1
          "1000000000001011" WHEN ADDR="00010100" AND CS_I='0' ELSE		--JNZ		JUDGE
          "1011001100000000" WHEN ADDR="00010101" AND CS_I='0' ELSE		--NEG		R3
          "1100110000000000" WHEN ADDR="00010110" AND CS_I='0' ELSE		--OUT		R3
          "0000000000000000";
END A;


